library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.constants_pkg.all;

entity rom_instr_test is
    clk : in std_logic
    write_address : out
