library ieee;
use ieee.std_logic_1164.all;

package constants_pkg is
    constant INSTR_MEM_LENGTH : integer := 5;
    constant DATA_LENGTH : integer := 64;
end package constants_pkg;

package body constants_pkg is
end package body constants_pkg;
