library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.constants_pkg.all;

entity top is
    port (

    );
end top;

architecture top_level of top is
-- component
 

begin



end top_level ; -- top